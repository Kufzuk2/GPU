module load_asm
#(
    parameter INSTR_SIZE = 16,
    parameter INSTR_NUM  = 288,
    parameter FULL_DEPTH = 1024
)
(
    input wire clk,
    input wire rst,

    output wire [INSTR_NUM * INSTR_SIZE - 1: 0] data_frames_line
);
    reg [INSTR_SIZE - 1: 0] data_frames [INSTR_NUM - 1: 0];
    

    genvar a;
    generate
        for (a = 0; a < INSTR_NUM; a = a + 1) begin : data_assign
            assign data_frames_line [INSTR_SIZE * (a + 1) - 1: INSTR_SIZE * a] = data_frames[a];
        end
    endgenerate


    always @(posedge clk) begin
        if (rst) begin
            data_frames[  0] <= 16'b0000000000000001;
            data_frames[  1] <= 16'b1111111111111110;
            data_frames[  2] <= 16'b1111111111111110;
            data_frames[  3] <= 16'b0000000000000000;
            data_frames[  4] <= 16'b0000000000000000;
            data_frames[  5] <= 16'b0000000000000000;
            data_frames[  6] <= 16'b0000000000000000;
            data_frames[  7] <= 16'b0000000000000000;
            data_frames[  8] <= 16'b0000000000000000;
            data_frames[  9] <= 16'b0000000000000000;
            data_frames[ 10] <= 16'b0000000000000000;
            data_frames[ 11] <= 16'b0000000000000000;
            data_frames[ 12] <= 16'b0000000000000000;
            data_frames[ 13] <= 16'b0000000000000000;
            data_frames[ 14] <= 16'b0000000000000000;
            data_frames[ 15] <= 16'b0000000000000000;
            data_frames[ 16] <= 16'b1100000000000011;
            data_frames[ 17] <= 16'b1100000001001001;
            data_frames[ 18] <= 16'b1100111111001010;
            data_frames[ 19] <= 16'b1100000000011100;
            data_frames[ 20] <= 16'b0000000000000000;
            data_frames[ 21] <= 16'b0000000000000000;
            data_frames[ 22] <= 16'b0000000000000000;
            data_frames[ 23] <= 16'b0000000000000000;
            data_frames[ 24] <= 16'b0000000000000000;
            data_frames[ 25] <= 16'b0000000000000000;
            data_frames[ 26] <= 16'b0000000000000000;
            data_frames[ 27] <= 16'b0000000000000000;
            data_frames[ 28] <= 16'b0000000000000000;
            data_frames[ 29] <= 16'b0000000000000000;
            data_frames[ 30] <= 16'b0000000000000000;
            data_frames[ 31] <= 16'b1111000000000000;
            data_frames[ 32] <= 16'b0000000000000001;
            data_frames[ 33] <= 16'b1111111111111110;
            data_frames[ 34] <= 16'b1111111111111110;
            data_frames[ 35] <= 16'b0000000000000000;
            data_frames[ 36] <= 16'b0000000000000000;
            data_frames[ 37] <= 16'b0000000000000000;
            data_frames[ 38] <= 16'b0000000000000000;
            data_frames[ 39] <= 16'b0000000000000000;
            data_frames[ 40] <= 16'b0000000000010000;
            data_frames[ 41] <= 16'b0010000000110000;
            data_frames[ 42] <= 16'b0100000001010000;
            data_frames[ 43] <= 16'b0110000001110000;
            data_frames[ 44] <= 16'b1000000010010000;
            data_frames[ 45] <= 16'b1010000010110000;
            data_frames[ 46] <= 16'b1100000011010000;
            data_frames[ 47] <= 16'b1110000011110000;
            data_frames[ 48] <= 16'b1101001111110000;
            data_frames[ 49] <= 16'b0001111111001111;
            data_frames[ 50] <= 16'b0011001110010110;
            data_frames[ 51] <= 16'b0010011011110100;
            data_frames[ 52] <= 16'b1110010000000000;
            data_frames[ 53] <= 16'b1101001111110000;
            data_frames[ 54] <= 16'b0001111111001111;
            data_frames[ 55] <= 16'b0001000010010000;
            data_frames[ 56] <= 16'b1101001111110000;
            data_frames[ 57] <= 16'b0001111111001111;
            data_frames[ 58] <= 16'b0010101000000100;
            data_frames[ 59] <= 16'b1110010001110000;
            data_frames[ 60] <= 16'b0000000000000000;
            data_frames[ 61] <= 16'b0000000000000000;
            data_frames[ 62] <= 16'b0000000000000000;
            data_frames[ 63] <= 16'b1111000000000000;
            data_frames[ 64] <= 16'b0000000000000001;
            data_frames[ 65] <= 16'b0000000000000001;
            data_frames[ 66] <= 16'b0000000000000001;
            data_frames[ 67] <= 16'b0000000000000000;
            data_frames[ 68] <= 16'b0000000000000000;
            data_frames[ 69] <= 16'b0000000000000000;
            data_frames[ 70] <= 16'b0000000000000000;
            data_frames[ 71] <= 16'b0000000000000000;
            data_frames[ 72] <= 16'b0000000000000000;
            data_frames[ 73] <= 16'b0000000000000000;
            data_frames[ 74] <= 16'b0000000000000000;
            data_frames[ 75] <= 16'b0000000000000000;
            data_frames[ 76] <= 16'b0000000000000000;
            data_frames[ 77] <= 16'b0000000000000000;
            data_frames[ 78] <= 16'b0000000000000000;
            data_frames[ 79] <= 16'b0000000000000000;
            data_frames[ 80] <= 16'b1100000000000011;
            data_frames[ 81] <= 16'b1100000001001001;
            data_frames[ 82] <= 16'b1100111111001010;
            data_frames[ 83] <= 16'b1100000000011100;
            data_frames[ 84] <= 16'b1101001111110000;
            data_frames[ 85] <= 16'b0001000010010000;
            data_frames[ 86] <= 16'b0001111111001111;
            data_frames[ 87] <= 16'b0010101000000100;
            data_frames[ 88] <= 16'b1110010001000000;
            data_frames[ 89] <= 16'b1101001111110000;
            data_frames[ 90] <= 16'b0001111111001111;
            data_frames[ 91] <= 16'b0001000010010000;
            data_frames[ 92] <= 16'b0000000000000000;
            data_frames[ 93] <= 16'b0000000000000000;
            data_frames[ 94] <= 16'b0000000000000000;
            data_frames[ 95] <= 16'b1111000000000000;
            data_frames[ 96] <= 16'b0000000000000001;
            data_frames[ 97] <= 16'b1111111111111111;
            data_frames[ 98] <= 16'b1111111111111111;
            data_frames[ 99] <= 16'b0000000000000000;
            data_frames[100] <= 16'b0000000000000000;
            data_frames[101] <= 16'b0000000000000000;
            data_frames[102] <= 16'b0000000000000000;
            data_frames[103] <= 16'b0000000000000000;
            data_frames[104] <= 16'b0000010000010100;
            data_frames[105] <= 16'b0010010000110100;
            data_frames[106] <= 16'b0100010001010100;
            data_frames[107] <= 16'b0110010001110100;
            data_frames[108] <= 16'b1000010010010100;
            data_frames[109] <= 16'b1010010010110100;
            data_frames[110] <= 16'b1100010011010100;
            data_frames[111] <= 16'b1110010011110100;
            data_frames[112] <= 16'b1100010000001000;
            data_frames[113] <= 16'b0011001110010101;
            data_frames[114] <= 16'b0001010111000101;
            data_frames[115] <= 16'b0001010110000101;
            data_frames[116] <= 16'b1101001111110000;
            data_frames[117] <= 16'b0001111111001111;
            data_frames[118] <= 16'b0010010111110100;
            data_frames[119] <= 16'b1110010001000000;
            data_frames[120] <= 16'b1101001111110000;
            data_frames[121] <= 16'b0001111111001111;
            data_frames[122] <= 16'b0001000010010000;
            data_frames[123] <= 16'b1101001111110000;
            data_frames[124] <= 16'b0001111111001111;
            data_frames[125] <= 16'b0010101000000100;
            data_frames[126] <= 16'b1110010010100000;
            data_frames[127] <= 16'b1111000000000000;
            data_frames[128] <= 16'b0000000000000001;
            data_frames[129] <= 16'b1111111111111111;
            data_frames[130] <= 16'b1111111111111111;
            data_frames[131] <= 16'b0000000000000000;
            data_frames[132] <= 16'b0000000000000000;
            data_frames[133] <= 16'b0000000000000000;
            data_frames[134] <= 16'b0000000000000000;
            data_frames[135] <= 16'b0000000000000000;
            data_frames[136] <= 16'b0000100000011000;
            data_frames[137] <= 16'b0010100000111000;
            data_frames[138] <= 16'b0100100001011000;
            data_frames[139] <= 16'b0110100001111000;
            data_frames[140] <= 16'b1000100010011000;
            data_frames[141] <= 16'b1010100010111000;
            data_frames[142] <= 16'b1100100011011000;
            data_frames[143] <= 16'b1110100011111000;
            data_frames[144] <= 16'b0001010111000101;
            data_frames[145] <= 16'b0001010110000101;
            data_frames[146] <= 16'b1101001111110000;
            data_frames[147] <= 16'b0001111111001111;
            data_frames[148] <= 16'b0010010111110100;
            data_frames[149] <= 16'b1110010000100000;
            data_frames[150] <= 16'b1101001111110000;
            data_frames[151] <= 16'b0001111111001111;
            data_frames[152] <= 16'b0001000010010000;
            data_frames[153] <= 16'b1101001111110000;
            data_frames[154] <= 16'b0001111111001111;
            data_frames[155] <= 16'b0010101000000100;
            data_frames[156] <= 16'b1110010010000000;
            data_frames[157] <= 16'b0000000000000000;
            data_frames[158] <= 16'b0000000000000000;
            data_frames[159] <= 16'b1111000000000000;
            data_frames[160] <= 16'b0000000000000001;
            data_frames[161] <= 16'b0111111111111111;
            data_frames[162] <= 16'b1111111111111111;
            data_frames[163] <= 16'b0000000000000000;
            data_frames[164] <= 16'b0000000000000000;
            data_frames[165] <= 16'b0000000000000000;
            data_frames[166] <= 16'b0000000000000000;
            data_frames[167] <= 16'b0000000000000000;
            data_frames[168] <= 16'b0000110000011100;
            data_frames[169] <= 16'b0010110000111100;
            data_frames[170] <= 16'b0100110001011100;
            data_frames[171] <= 16'b0110110001111100;
            data_frames[172] <= 16'b1000110010011100;
            data_frames[173] <= 16'b1010110010111100;
            data_frames[174] <= 16'b1100110011011100;
            data_frames[175] <= 16'b1110110011111100;
            data_frames[176] <= 16'b0001010111000101;
            data_frames[177] <= 16'b0001010110000101;
            data_frames[178] <= 16'b1101001111110000;
            data_frames[179] <= 16'b0001111111001111;
            data_frames[180] <= 16'b0010010111110100;
            data_frames[181] <= 16'b1110010000100000;
            data_frames[182] <= 16'b1101001111110000;
            data_frames[183] <= 16'b0001111111001111;
            data_frames[184] <= 16'b0001000010010000;
            data_frames[185] <= 16'b1101001111110000;
            data_frames[186] <= 16'b0001111111001111;
            data_frames[187] <= 16'b0010101000000100;
            data_frames[188] <= 16'b1110010010000000;
            data_frames[189] <= 16'b0000000000000000;
            data_frames[190] <= 16'b0000000000000000;
            data_frames[191] <= 16'b1111000000000000;
            data_frames[192] <= 16'b0000000000000001;
            data_frames[193] <= 16'b1000000000000000;
            data_frames[194] <= 16'b1000000000000000;
            data_frames[195] <= 16'b0000000000000000;
            data_frames[196] <= 16'b0000000000000000;
            data_frames[197] <= 16'b0000000000000000;
            data_frames[198] <= 16'b0000000000000000;
            data_frames[199] <= 16'b0000000000000000;
            data_frames[200] <= 16'b0000000000000000;
            data_frames[201] <= 16'b0000000000000000;
            data_frames[202] <= 16'b0000000000000000;
            data_frames[203] <= 16'b0000000000000000;
            data_frames[204] <= 16'b0000000000000000;
            data_frames[205] <= 16'b0000000000000000;
            data_frames[206] <= 16'b0000000000000000;
            data_frames[207] <= 16'b0000000000000000;
            data_frames[208] <= 16'b0001010111000101;
            data_frames[209] <= 16'b0001010110000101;
            data_frames[210] <= 16'b1101001111111010;
            data_frames[211] <= 16'b0001111111001111;
            data_frames[212] <= 16'b0010010111110100;
            data_frames[213] <= 16'b1110010000100000;
            data_frames[214] <= 16'b1101001111111010;
            data_frames[215] <= 16'b0000000000000000;
            data_frames[216] <= 16'b0000000000000000;
            data_frames[217] <= 16'b0000000000000000;
            data_frames[218] <= 16'b0000000000000000;
            data_frames[219] <= 16'b0000000000000000;
            data_frames[220] <= 16'b0000000000000000;
            data_frames[221] <= 16'b0000000000000000;
            data_frames[222] <= 16'b0000000000000000;
            data_frames[223] <= 16'b1111000000000000;
            data_frames[224] <= 16'b0000000000000001;
            data_frames[225] <= 16'b1111111111111111;
            data_frames[226] <= 16'b1111111111111111;
            data_frames[227] <= 16'b0000000000000000;
            data_frames[228] <= 16'b0000000000000000;
            data_frames[229] <= 16'b0000000000000000;
            data_frames[230] <= 16'b0000000000000000;
            data_frames[231] <= 16'b0000000000000000;
            data_frames[232] <= 16'b0000000000000000;
            data_frames[233] <= 16'b0000000000000000;
            data_frames[234] <= 16'b0000000000000000;
            data_frames[235] <= 16'b0000000000000000;
            data_frames[236] <= 16'b0000000000000000;
            data_frames[237] <= 16'b0000000000000000;
            data_frames[238] <= 16'b0000000000000000;
            data_frames[239] <= 16'b0000000000000000;
            data_frames[240] <= 16'b1100000000000011;
            data_frames[241] <= 16'b1100000001001001;
            data_frames[242] <= 16'b1100111111111010;
            data_frames[243] <= 16'b1100000000011100;
            data_frames[244] <= 16'b1100000000001011;
            data_frames[245] <= 16'b1100000000001111;
            data_frames[246] <= 16'b0000000000000000;
            data_frames[247] <= 16'b0000000000000000;
            data_frames[248] <= 16'b0000000000000000;
            data_frames[249] <= 16'b0000000000000000;
            data_frames[250] <= 16'b0000000000000000;
            data_frames[251] <= 16'b0000000000000000;
            data_frames[252] <= 16'b0000000000000000;
            data_frames[253] <= 16'b0000000000000000;
            data_frames[254] <= 16'b0000000000000000;
            data_frames[255] <= 16'b1111000000000000;
            data_frames[256] <= 16'b0000000000000001;
            data_frames[257] <= 16'b1111111111111111;
            data_frames[258] <= 16'b1111111111111111;
            data_frames[259] <= 16'b0000000000000000;
            data_frames[260] <= 16'b0000000000000000;
            data_frames[261] <= 16'b0000000000000000;
            data_frames[262] <= 16'b0000000000000000;
            data_frames[263] <= 16'b0000000000000000;
            data_frames[264] <= 16'b0000000000000000;
            data_frames[265] <= 16'b0000000000000000;
            data_frames[266] <= 16'b0000000000000000;
            data_frames[267] <= 16'b0000000000000000;
            data_frames[268] <= 16'b0000000000000000;
            data_frames[269] <= 16'b0000000000000000;
            data_frames[270] <= 16'b0000000000000000;
            data_frames[271] <= 16'b0000000000000000;
            data_frames[272] <= 16'b0000000000000000;
            data_frames[273] <= 16'b1011001111110101;
            data_frames[274] <= 16'b0001010110010110;
            data_frames[275] <= 16'b1101001111110110;
            data_frames[276] <= 16'b0001111111001111;
            data_frames[277] <= 16'b0010101011111000;
            data_frames[278] <= 16'b1110100000010000;
            data_frames[279] <= 16'b1011001111110101;
            data_frames[280] <= 16'b0001010110010110;
            data_frames[281] <= 16'b1101001111110110;
            data_frames[282] <= 16'b0000000000000000;
            data_frames[283] <= 16'b0000000000000000;
            data_frames[284] <= 16'b0000000000000000;
            data_frames[285] <= 16'b0000000000000000;
            data_frames[286] <= 16'b0000000000000000;
            data_frames[287] <= 16'b1111000000000000;
        end else begin
            data_frames[  0] <= data_frames[  0];
            data_frames[  1] <= data_frames[  1];
            data_frames[  2] <= data_frames[  2];
            data_frames[  3] <= data_frames[  3];
            data_frames[  4] <= data_frames[  4];
            data_frames[  5] <= data_frames[  5];
            data_frames[  6] <= data_frames[  6];
            data_frames[  7] <= data_frames[  7];
            data_frames[  8] <= data_frames[  8];
            data_frames[  9] <= data_frames[  9];
            data_frames[ 10] <= data_frames[ 10];
            data_frames[ 11] <= data_frames[ 11];
            data_frames[ 12] <= data_frames[ 12];
            data_frames[ 13] <= data_frames[ 13];
            data_frames[ 14] <= data_frames[ 14];
            data_frames[ 15] <= data_frames[ 15];
            data_frames[ 16] <= data_frames[ 16];
            data_frames[ 17] <= data_frames[ 17];
            data_frames[ 18] <= data_frames[ 18];
            data_frames[ 19] <= data_frames[ 19];
            data_frames[ 20] <= data_frames[ 20];
            data_frames[ 21] <= data_frames[ 21];
            data_frames[ 22] <= data_frames[ 22];
            data_frames[ 23] <= data_frames[ 23];
            data_frames[ 24] <= data_frames[ 24];
            data_frames[ 25] <= data_frames[ 25];
            data_frames[ 26] <= data_frames[ 26];
            data_frames[ 27] <= data_frames[ 27];
            data_frames[ 28] <= data_frames[ 28];
            data_frames[ 29] <= data_frames[ 29];
            data_frames[ 30] <= data_frames[ 30];
            data_frames[ 31] <= data_frames[ 31];
            data_frames[ 32] <= data_frames[ 32];
            data_frames[ 33] <= data_frames[ 33];
            data_frames[ 34] <= data_frames[ 34];
            data_frames[ 35] <= data_frames[ 35];
            data_frames[ 36] <= data_frames[ 36];
            data_frames[ 37] <= data_frames[ 37];
            data_frames[ 38] <= data_frames[ 38];
            data_frames[ 39] <= data_frames[ 39];
            data_frames[ 40] <= data_frames[ 40];
            data_frames[ 41] <= data_frames[ 41];
            data_frames[ 42] <= data_frames[ 42];
            data_frames[ 43] <= data_frames[ 43];
            data_frames[ 44] <= data_frames[ 44];
            data_frames[ 45] <= data_frames[ 45];
            data_frames[ 46] <= data_frames[ 46];
            data_frames[ 47] <= data_frames[ 47];
            data_frames[ 48] <= data_frames[ 48];
            data_frames[ 49] <= data_frames[ 49];
            data_frames[ 50] <= data_frames[ 50];
            data_frames[ 51] <= data_frames[ 51];
            data_frames[ 52] <= data_frames[ 52];
            data_frames[ 53] <= data_frames[ 53];
            data_frames[ 54] <= data_frames[ 54];
            data_frames[ 55] <= data_frames[ 55];
            data_frames[ 56] <= data_frames[ 56];
            data_frames[ 57] <= data_frames[ 57];
            data_frames[ 58] <= data_frames[ 58];
            data_frames[ 59] <= data_frames[ 59];
            data_frames[ 60] <= data_frames[ 60];
            data_frames[ 61] <= data_frames[ 61];
            data_frames[ 62] <= data_frames[ 62];
            data_frames[ 63] <= data_frames[ 63];
            data_frames[ 64] <= data_frames[ 64];
            data_frames[ 65] <= data_frames[ 65];
            data_frames[ 66] <= data_frames[ 66];
            data_frames[ 67] <= data_frames[ 67];
            data_frames[ 68] <= data_frames[ 68];
            data_frames[ 69] <= data_frames[ 69];
            data_frames[ 70] <= data_frames[ 70];
            data_frames[ 71] <= data_frames[ 71];
            data_frames[ 72] <= data_frames[ 72];
            data_frames[ 73] <= data_frames[ 73];
            data_frames[ 74] <= data_frames[ 74];
            data_frames[ 75] <= data_frames[ 75];
            data_frames[ 76] <= data_frames[ 76];
            data_frames[ 77] <= data_frames[ 77];
            data_frames[ 78] <= data_frames[ 78];
            data_frames[ 79] <= data_frames[ 79];
            data_frames[ 80] <= data_frames[ 80];
            data_frames[ 81] <= data_frames[ 81];
            data_frames[ 82] <= data_frames[ 82];
            data_frames[ 83] <= data_frames[ 83];
            data_frames[ 84] <= data_frames[ 84];
            data_frames[ 85] <= data_frames[ 85];
            data_frames[ 86] <= data_frames[ 86];
            data_frames[ 87] <= data_frames[ 87];
            data_frames[ 88] <= data_frames[ 88];
            data_frames[ 89] <= data_frames[ 89];
            data_frames[ 90] <= data_frames[ 90];
            data_frames[ 91] <= data_frames[ 91];
            data_frames[ 92] <= data_frames[ 92];
            data_frames[ 93] <= data_frames[ 93];
            data_frames[ 94] <= data_frames[ 94];
            data_frames[ 95] <= data_frames[ 95];
            data_frames[ 96] <= data_frames[ 96];
            data_frames[ 97] <= data_frames[ 97];
            data_frames[ 98] <= data_frames[ 98];
            data_frames[ 99] <= data_frames[ 99];
            data_frames[100] <= data_frames[100];
            data_frames[101] <= data_frames[101];
            data_frames[102] <= data_frames[102];
            data_frames[103] <= data_frames[103];
            data_frames[104] <= data_frames[104];
            data_frames[105] <= data_frames[105];
            data_frames[106] <= data_frames[106];
            data_frames[107] <= data_frames[107];
            data_frames[108] <= data_frames[108];
            data_frames[109] <= data_frames[109];
            data_frames[110] <= data_frames[110];
            data_frames[111] <= data_frames[111];
            data_frames[112] <= data_frames[112];
            data_frames[113] <= data_frames[113];
            data_frames[114] <= data_frames[114];
            data_frames[115] <= data_frames[115];
            data_frames[116] <= data_frames[116];
            data_frames[117] <= data_frames[117];
            data_frames[118] <= data_frames[118];
            data_frames[119] <= data_frames[119];
            data_frames[120] <= data_frames[120];
            data_frames[121] <= data_frames[121];
            data_frames[122] <= data_frames[122];
            data_frames[123] <= data_frames[123];
            data_frames[124] <= data_frames[124];
            data_frames[125] <= data_frames[125];
            data_frames[126] <= data_frames[126];
            data_frames[127] <= data_frames[127];
            data_frames[128] <= data_frames[128];
            data_frames[129] <= data_frames[129];
            data_frames[130] <= data_frames[130];
            data_frames[131] <= data_frames[131];
            data_frames[132] <= data_frames[132];
            data_frames[133] <= data_frames[133];
            data_frames[134] <= data_frames[134];
            data_frames[135] <= data_frames[135];
            data_frames[136] <= data_frames[136];
            data_frames[137] <= data_frames[137];
            data_frames[138] <= data_frames[138];
            data_frames[139] <= data_frames[139];
            data_frames[140] <= data_frames[140];
            data_frames[141] <= data_frames[141];
            data_frames[142] <= data_frames[142];
            data_frames[143] <= data_frames[143];
            data_frames[144] <= data_frames[144];
            data_frames[145] <= data_frames[145];
            data_frames[146] <= data_frames[146];
            data_frames[147] <= data_frames[147];
            data_frames[148] <= data_frames[148];
            data_frames[149] <= data_frames[149];
            data_frames[150] <= data_frames[150];
            data_frames[151] <= data_frames[151];
            data_frames[152] <= data_frames[152];
            data_frames[153] <= data_frames[153];
            data_frames[154] <= data_frames[154];
            data_frames[155] <= data_frames[155];
            data_frames[156] <= data_frames[156];
            data_frames[157] <= data_frames[157];
            data_frames[158] <= data_frames[158];
            data_frames[159] <= data_frames[159];
            data_frames[160] <= data_frames[160];
            data_frames[161] <= data_frames[161];
            data_frames[162] <= data_frames[162];
            data_frames[163] <= data_frames[163];
            data_frames[164] <= data_frames[164];
            data_frames[165] <= data_frames[165];
            data_frames[166] <= data_frames[166];
            data_frames[167] <= data_frames[167];
            data_frames[168] <= data_frames[168];
            data_frames[169] <= data_frames[169];
            data_frames[170] <= data_frames[170];
            data_frames[171] <= data_frames[171];
            data_frames[172] <= data_frames[172];
            data_frames[173] <= data_frames[173];
            data_frames[174] <= data_frames[174];
            data_frames[175] <= data_frames[175];
            data_frames[176] <= data_frames[176];
            data_frames[177] <= data_frames[177];
            data_frames[178] <= data_frames[178];
            data_frames[179] <= data_frames[179];
            data_frames[180] <= data_frames[180];
            data_frames[181] <= data_frames[181];
            data_frames[182] <= data_frames[182];
            data_frames[183] <= data_frames[183];
            data_frames[184] <= data_frames[184];
            data_frames[185] <= data_frames[185];
            data_frames[186] <= data_frames[186];
            data_frames[187] <= data_frames[187];
            data_frames[188] <= data_frames[188];
            data_frames[189] <= data_frames[189];
            data_frames[190] <= data_frames[190];
            data_frames[191] <= data_frames[191];
            data_frames[192] <= data_frames[192];
            data_frames[193] <= data_frames[193];
            data_frames[194] <= data_frames[194];
            data_frames[195] <= data_frames[195];
            data_frames[196] <= data_frames[196];
            data_frames[197] <= data_frames[197];
            data_frames[198] <= data_frames[198];
            data_frames[199] <= data_frames[199];
            data_frames[200] <= data_frames[200];
            data_frames[201] <= data_frames[201];
            data_frames[202] <= data_frames[202];
            data_frames[203] <= data_frames[203];
            data_frames[204] <= data_frames[204];
            data_frames[205] <= data_frames[205];
            data_frames[206] <= data_frames[206];
            data_frames[207] <= data_frames[207];
            data_frames[208] <= data_frames[208];
            data_frames[209] <= data_frames[209];
            data_frames[210] <= data_frames[210];
            data_frames[211] <= data_frames[211];
            data_frames[212] <= data_frames[212];
            data_frames[213] <= data_frames[213];
            data_frames[214] <= data_frames[214];
            data_frames[215] <= data_frames[215];
            data_frames[216] <= data_frames[216];
            data_frames[217] <= data_frames[217];
            data_frames[218] <= data_frames[218];
            data_frames[219] <= data_frames[219];
            data_frames[220] <= data_frames[220];
            data_frames[221] <= data_frames[221];
            data_frames[222] <= data_frames[222];
            data_frames[223] <= data_frames[223];
            data_frames[224] <= data_frames[224];
            data_frames[225] <= data_frames[225];
            data_frames[226] <= data_frames[226];
            data_frames[227] <= data_frames[227];
            data_frames[228] <= data_frames[228];
            data_frames[229] <= data_frames[229];
            data_frames[230] <= data_frames[230];
            data_frames[231] <= data_frames[231];
            data_frames[232] <= data_frames[232];
            data_frames[233] <= data_frames[233];
            data_frames[234] <= data_frames[234];
            data_frames[235] <= data_frames[235];
            data_frames[236] <= data_frames[236];
            data_frames[237] <= data_frames[237];
            data_frames[238] <= data_frames[238];
            data_frames[239] <= data_frames[239];
            data_frames[240] <= data_frames[240];
            data_frames[241] <= data_frames[241];
            data_frames[242] <= data_frames[242];
            data_frames[243] <= data_frames[243];
            data_frames[244] <= data_frames[244];
            data_frames[245] <= data_frames[245];
            data_frames[246] <= data_frames[246];
            data_frames[247] <= data_frames[247];
            data_frames[248] <= data_frames[248];
            data_frames[249] <= data_frames[249];
            data_frames[250] <= data_frames[250];
            data_frames[251] <= data_frames[251];
            data_frames[252] <= data_frames[252];
            data_frames[253] <= data_frames[253];
            data_frames[254] <= data_frames[254];
            data_frames[255] <= data_frames[255];
            data_frames[256] <= data_frames[256];
            data_frames[257] <= data_frames[257];
            data_frames[258] <= data_frames[258];
            data_frames[259] <= data_frames[259];
            data_frames[260] <= data_frames[260];
            data_frames[261] <= data_frames[261];
            data_frames[262] <= data_frames[262];
            data_frames[263] <= data_frames[263];
            data_frames[264] <= data_frames[264];
            data_frames[265] <= data_frames[265];
            data_frames[266] <= data_frames[266];
            data_frames[267] <= data_frames[267];
            data_frames[268] <= data_frames[268];
            data_frames[269] <= data_frames[269];
            data_frames[270] <= data_frames[270];
            data_frames[271] <= data_frames[271];
            data_frames[272] <= data_frames[272];
            data_frames[273] <= data_frames[273];
            data_frames[274] <= data_frames[274];
            data_frames[275] <= data_frames[275];
            data_frames[276] <= data_frames[276];
            data_frames[277] <= data_frames[277];
            data_frames[278] <= data_frames[278];
            data_frames[279] <= data_frames[279];
            data_frames[280] <= data_frames[280];
            data_frames[281] <= data_frames[281];
            data_frames[282] <= data_frames[282];
            data_frames[283] <= data_frames[283];
            data_frames[284] <= data_frames[284];
            data_frames[285] <= data_frames[285];
            data_frames[286] <= data_frames[286];
            data_frames[287] <= data_frames[287];
        end
    end

endmodule
